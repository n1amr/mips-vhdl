library IEEE;
use IEEE.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_textio.all;
use std.textio.all;

entity DataMemory is
  port( address : in std_logic_vector(31 downto 0);
        clk : in std_logic ;
        write_data: in std_logic_vector(31 downto 0);
        MemWrite, MemRead: in std_logic;
        read_data : out std_logic_vector(31 downto 0)
      );
end entity;

architecture bev of DataMemory is
  type memory is array (0 to 255) of std_logic_vector(7 downto 0);
  signal mem : memory;
begin
  process(clk)
  begin
    if(clk'event and clk = '1' and MemWrite = '1') then
      mem(conv_integer(address)) <= write_data(31 downto 24);
      mem(conv_integer(address) + 1) <= write_data(23 downto 16);
      mem(conv_integer(address) + 2) <= write_data(15 downto 8);
      mem(conv_integer(address) + 3) <= write_data(7 downto 0);
    end if;
  end process;
  
  process(MemRead, address)
  begin
    if(MemRead = '1') then
      read_data(31 downto 24) <= mem(conv_integer(address));
      read_data(23 downto 16) <= mem(conv_integer(address) + 1);
      read_data(15 downto 8) <= mem(conv_integer(address) + 2);
      read_data(7 downto 0) <= mem(conv_integer(address) + 3);
    end if;
  end process;

  --process
  --  constant FILENAME : string :="data-memory.mem";
  --  FILE mFile : TEXT;
  --  variable i : integer := 0;
  --  variable mLIne : LINE;
  --  variable mByte : std_logic_vector(7 downto 0);
  --begin
  --  File_Open(mFile, FILENAME, read_mode);
  --  while( (i <= 15) and (not EndFile(mFile))) loop
  --    readline (mFile, mLIne);
  --    next when mLIne(1) = '#';
  --    read(mLIne, mByte);
  --    mem(i) <= mByte;
  --    i := i + 1;
  --  end loop;
    
  --  File_Close(mFile);
  --  wait;
  --end process;
end bev;
