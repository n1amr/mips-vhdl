library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
entity adder is
  port (  a : in bit_vector (31 DOWNTO 0);
          b : in bit_vector (31 DOWNTO 0);
          result : out bit_vector (31 DOWNTO 0));
end adder;

architecture behave of adder is
begin
  result <= a + b;
end behave;

